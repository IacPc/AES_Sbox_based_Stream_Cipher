module sbox_lut(lut_in);
	input  [7:0] lut_in;
	output [7:0] lut_out;

	always @(lut_in) begin
		case (lut_in)
			8'h00: lut_out <= 8'h63; 
			8'h01: lut_out <= 8'h7c; 
			8'h02: lut_out <= 8'h77; 
			8'h03: lut_out <= 8'h7b; 
			8'h04: lut_out <= 8'hf2; 
			8'h05: lut_out <= 8'h6b; 
			8'h06: lut_out <= 8'h6f; 
			8'h07: lut_out <= 8'hc5; 
			8'h08: lut_out <= 8'h30; 
			8'h09: lut_out <= 8'h01; 
			8'h0a: lut_out <= 8'h67; 
			8'h0b: lut_out <= 8'h2b; 
			8'h0c: lut_out <= 8'hfe; 
			8'h0d: lut_out <= 8'hd7; 
			8'h0e: lut_out <= 8'hab; 
			8'h0f: lut_out <= 8'h76; 
			8'h10: lut_out <= 8'hca; 
			8'h11: lut_out <= 8'h82; 
			8'h12: lut_out <= 8'hc9; 
			8'h13: lut_out <= 8'h7d; 
			8'h14: lut_out <= 8'hfa; 
			8'h15: lut_out <= 8'h59; 
			8'h16: lut_out <= 8'h47; 
			8'h17: lut_out <= 8'hf0; 
			8'h18: lut_out <= 8'had; 
			8'h19: lut_out <= 8'hd4; 
			8'h1a: lut_out <= 8'ha2; 
			8'h1b: lut_out <= 8'haf; 
			8'h1c: lut_out <= 8'h9c; 
			8'h1d: lut_out <= 8'ha4; 
			8'h1e: lut_out <= 8'h72; 
			8'h1f: lut_out <= 8'hc0; 
			8'h20: lut_out <= 8'hb7; 
			8'h21: lut_out <= 8'hfd; 
			8'h22: lut_out <= 8'h93; 
			8'h23: lut_out <= 8'h26; 
			8'h24: lut_out <= 8'h36; 
			8'h25: lut_out <= 8'h3f; 
			8'h26: lut_out <= 8'hf7; 
			8'h27: lut_out <= 8'hcc; 
			8'h28: lut_out <= 8'h34; 
			8'h29: lut_out <= 8'ha5; 
			8'h2a: lut_out <= 8'he5; 
			8'h2b: lut_out <= 8'hf1; 
			8'h2c: lut_out <= 8'h71; 
			8'h2d: lut_out <= 8'hd8; 
			8'h2e: lut_out <= 8'h31; 
			8'h2f: lut_out <= 8'h15; 
			8'h30: lut_out <= 8'h04; 
			8'h31: lut_out <= 8'hc7; 
			8'h32: lut_out <= 8'h23; 
			8'h33: lut_out <= 8'hc3; 
			8'h34: lut_out <= 8'h18; 
			8'h35: lut_out <= 8'h96; 
			8'h36: lut_out <= 8'h05; 
			8'h37: lut_out <= 8'h9a; 
			8'h38: lut_out <= 8'h07; 
			8'h39: lut_out <= 8'h12; 
			8'h3a: lut_out <= 8'h80; 
			8'h3b: lut_out <= 8'he2; 
			8'h3c: lut_out <= 8'heb; 
			8'h3d: lut_out <= 8'h27; 
			8'h3e: lut_out <= 8'hb2; 
			8'h3f: lut_out <= 8'h75; 
			8'h40: lut_out <= 8'h09; 
			8'h41: lut_out <= 8'h83; 
			8'h42: lut_out <= 8'h2c; 
			8'h43: lut_out <= 8'h1a; 
			8'h44: lut_out <= 8'h1b; 
			8'h45: lut_out <= 8'h6e; 
			8'h46: lut_out <= 8'h5a; 
			8'h47: lut_out <= 8'ha0; 
			8'h48: lut_out <= 8'h52; 
			8'h49: lut_out <= 8'h3b; 
			8'h4a: lut_out <= 8'hd6; 
			8'h4b: lut_out <= 8'hb3; 
			8'h4c: lut_out <= 8'h29; 
			8'h4d: lut_out <= 8'he3; 
			8'h4e: lut_out <= 8'h2f; 
			8'h4f: lut_out <= 8'h84; 
			8'h50: lut_out <= 8'h53; 
			8'h51: lut_out <= 8'hd1; 
			8'h52: lut_out <= 8'h00; 
			8'h53: lut_out <= 8'hed; 
			8'h54: lut_out <= 8'h20; 
			8'h55: lut_out <= 8'hfc; 
			8'h56: lut_out <= 8'hb1; 
			8'h57: lut_out <= 8'h5b; 
			8'h58: lut_out <= 8'h6a; 
			8'h59: lut_out <= 8'hcb; 
			8'h5a: lut_out <= 8'hbe; 
			8'h5b: lut_out <= 8'h39; 
			8'h5c: lut_out <= 8'h4a; 
			8'h5d: lut_out <= 8'h4c; 
			8'h5e: lut_out <= 8'h58; 
			8'h5f: lut_out <= 8'hcf; 
			8'h60: lut_out <= 8'hd0; 
			8'h61: lut_out <= 8'hef; 
			8'h62: lut_out <= 8'haa; 
			8'h63: lut_out <= 8'hfb; 
			8'h64: lut_out <= 8'h43; 
			8'h65: lut_out <= 8'h4d; 
			8'h66: lut_out <= 8'h33; 
			8'h67: lut_out <= 8'h85; 
			8'h68: lut_out <= 8'h45; 
			8'h69: lut_out <= 8'hf9; 
			8'h6a: lut_out <= 8'h02; 
			8'h6b: lut_out <= 8'h7f; 
			8'h6c: lut_out <= 8'h50; 
			8'h6d: lut_out <= 8'h3c; 
			8'h6e: lut_out <= 8'h9f; 
			8'h6f: lut_out <= 8'ha8; 
			8'h70: lut_out <= 8'h51; 
			8'h71: lut_out <= 8'ha3; 
			8'h72: lut_out <= 8'h40; 
			8'h73: lut_out <= 8'h8f; 
			8'h74: lut_out <= 8'h92; 
			8'h75: lut_out <= 8'h9d; 
			8'h76: lut_out <= 8'h38; 
			8'h77: lut_out <= 8'hf5; 
			8'h78: lut_out <= 8'hbc; 
			8'h79: lut_out <= 8'hb6; 
			8'h7a: lut_out <= 8'hda; 
			8'h7b: lut_out <= 8'h21; 
			8'h7c: lut_out <= 8'h10; 
			8'h7d: lut_out <= 8'hff; 
			8'h7e: lut_out <= 8'hf3; 
			8'h7f: lut_out <= 8'hd2; 
			8'h80: lut_out <= 8'hcd; 
			8'h81: lut_out <= 8'h0c; 
			8'h82: lut_out <= 8'h13; 
			8'h83: lut_out <= 8'hec; 
			8'h84: lut_out <= 8'h5f; 
			8'h85: lut_out <= 8'h97; 
			8'h86: lut_out <= 8'h44; 
			8'h87: lut_out <= 8'h17; 
			8'h88: lut_out <= 8'hc4; 
			8'h89: lut_out <= 8'ha7; 
			8'h8a: lut_out <= 8'h7e; 
			8'h8b: lut_out <= 8'h3d; 
			8'h8c: lut_out <= 8'h64; 
			8'h8d: lut_out <= 8'h5d; 
			8'h8e: lut_out <= 8'h19; 
			8'h8f: lut_out <= 8'h73; 
			8'h90: lut_out <= 8'h60; 
			8'h91: lut_out <= 8'h81; 
			8'h92: lut_out <= 8'h4f; 
			8'h93: lut_out <= 8'hdc; 
			8'h94: lut_out <= 8'h22; 
			8'h95: lut_out <= 8'h2a; 
			8'h96: lut_out <= 8'h90; 
			8'h97: lut_out <= 8'h88; 
			8'h98: lut_out <= 8'h46; 
			8'h99: lut_out <= 8'hee; 
			8'h9a: lut_out <= 8'hb8; 
			8'h9b: lut_out <= 8'h14; 
			8'h9c: lut_out <= 8'hde; 
			8'h9d: lut_out <= 8'h5e; 
			8'h9e: lut_out <= 8'h0b; 
			8'h9f: lut_out <= 8'hdb; 
			8'ha0: lut_out <= 8'he0; 
			8'ha1: lut_out <= 8'h32; 
			8'ha2: lut_out <= 8'h3a; 
			8'ha3: lut_out <= 8'h0a; 
			8'ha4: lut_out <= 8'h49; 
			8'ha5: lut_out <= 8'h06; 
			8'ha6: lut_out <= 8'h24; 
			8'ha7: lut_out <= 8'h5c; 
			8'ha8: lut_out <= 8'hc2; 
			8'ha9: lut_out <= 8'hd3; 
			8'haa: lut_out <= 8'hac; 
			8'hab: lut_out <= 8'h62; 
			8'hac: lut_out <= 8'h91; 
			8'had: lut_out <= 8'h95; 
			8'hae: lut_out <= 8'he4; 
			8'haf: lut_out <= 8'h79; 
			8'hb0: lut_out <= 8'he7; 
			8'hb1: lut_out <= 8'hc8; 
			8'hb2: lut_out <= 8'h37; 
			8'hb3: lut_out <= 8'h6d; 
			8'hb4: lut_out <= 8'h8d; 
			8'hb5: lut_out <= 8'hd5; 
			8'hb6: lut_out <= 8'h4e; 
			8'hb7: lut_out <= 8'ha9; 
			8'hb8: lut_out <= 8'h6c; 
			8'hb9: lut_out <= 8'h56; 
			8'hba: lut_out <= 8'hf4; 
			8'hbb: lut_out <= 8'hea; 
			8'hbc: lut_out <= 8'h65; 
			8'hbd: lut_out <= 8'h7a; 
			8'hbe: lut_out <= 8'hae; 
			8'hbf: lut_out <= 8'h08; 
			8'hc0: lut_out <= 8'hba; 
			8'hc1: lut_out <= 8'h78; 
			8'hc2: lut_out <= 8'h25; 
			8'hc3: lut_out <= 8'h2e; 
			8'hc4: lut_out <= 8'h1c; 
			8'hc5: lut_out <= 8'ha6; 
			8'hc6: lut_out <= 8'hb4; 
			8'hc7: lut_out <= 8'hc6; 
			8'hc8: lut_out <= 8'he8; 
			8'hc9: lut_out <= 8'hdd; 
			8'hca: lut_out <= 8'h74; 
			8'hcb: lut_out <= 8'h1f; 
			8'hcc: lut_out <= 8'h4b; 
			8'hcd: lut_out <= 8'hbd; 
			8'hce: lut_out <= 8'h8b; 
			8'hcf: lut_out <= 8'h8a; 
			8'hd0: lut_out <= 8'h70; 
			8'hd1: lut_out <= 8'h3e; 
			8'hd2: lut_out <= 8'hb5; 
			8'hd3: lut_out <= 8'h66; 
			8'hd4: lut_out <= 8'h48; 
			8'hd5: lut_out <= 8'h03; 
			8'hd6: lut_out <= 8'hf6; 
			8'hd7: lut_out <= 8'h0e; 
			8'hd8: lut_out <= 8'h61; 
			8'hd9: lut_out <= 8'h35; 
			8'hda: lut_out <= 8'h57; 
			8'hdb: lut_out <= 8'hb9; 
			8'hdc: lut_out <= 8'h86; 
			8'hdd: lut_out <= 8'hc1; 
			8'hde: lut_out <= 8'h1d; 
			8'hdf: lut_out <= 8'h9e; 
			8'he0: lut_out <= 8'he1; 
			8'he1: lut_out <= 8'hf8; 
			8'he2: lut_out <= 8'h98; 
			8'he3: lut_out <= 8'h11; 
			8'he4: lut_out <= 8'h69; 
			8'he5: lut_out <= 8'hd9; 
			8'he6: lut_out <= 8'h8e; 
			8'he7: lut_out <= 8'h94; 
			8'he8: lut_out <= 8'h9b; 
			8'he9: lut_out <= 8'h1e; 
			8'hea: lut_out <= 8'h87; 
			8'heb: lut_out <= 8'he9; 
			8'hec: lut_out <= 8'hce; 
			8'hed: lut_out <= 8'h55; 
			8'hee: lut_out <= 8'h28; 
			8'hef: lut_out <= 8'hdf; 
			8'hf0: lut_out <= 8'h8c; 
			8'hf1: lut_out <= 8'ha1; 
			8'hf2: lut_out <= 8'h89; 
			8'hf3: lut_out <= 8'h0d; 
			8'hf4: lut_out <= 8'hbf; 
			8'hf5: lut_out <= 8'he6; 
			8'hf6: lut_out <= 8'h42; 
			8'hf7: lut_out <= 8'h68; 
			8'hf8: lut_out <= 8'h41; 
			8'hf9: lut_out <= 8'h99; 
			8'hfa: lut_out <= 8'h2d; 
			8'hfb: lut_out <= 8'h0f; 
			8'hfc: lut_out <= 8'hb0; 
			8'hfd: lut_out <= 8'h54; 
			8'hfe: lut_out <= 8'hbb; 
			8'hff: lut_out <= 8'h16; 
		endcase
	end
endmodule
